library verilog;
use verilog.vl_types.all;
entity Projeto_final_vlg_vec_tst is
end Projeto_final_vlg_vec_tst;
